* /home/roshan/eSim-Workspace/calc16/calc16.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Jul  2 17:30:09 2023

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ calcu16		
v1  clk GND pulse		
U2  clk Net-_U1-Pad1_ adc_bridge_1		
U3  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ 1 2 3 4 5 6 7 8 dac_bridge_8		
U4  Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ 9 10 11 12 13 14 15 16 dac_bridge_8		
U5  1 plot_v1		
U6  2 plot_v1		
U7  3 plot_v1		
U8  4 plot_v1		
U9  5 plot_v1		
U10  6 plot_v1		
U11  7 plot_v1		
U12  8 plot_v1		
U13  9 plot_v1		
U14  10 plot_v1		
U15  11 plot_v1		
U16  12 plot_v1		
U17  13 plot_v1		
U18  14 plot_v1		
U19  15 plot_v1		
U20  16 plot_v1		

.end
